library verilog;
use verilog.vl_types.all;
entity Test is
end Test;
