library verilog;
use verilog.vl_types.all;
entity FIR_TB is
end FIR_TB;
