library verilog;
use verilog.vl_types.all;
entity cordic_10_tb is
end cordic_10_tb;
