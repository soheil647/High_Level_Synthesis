library verilog;
use verilog.vl_types.all;
entity cordic_tb is
end cordic_tb;
