library verilog;
use verilog.vl_types.all;
entity Tseries_tb is
end Tseries_tb;
