library verilog;
use verilog.vl_types.all;
entity Absulote_tb is
end Absulote_tb;
