library verilog;
use verilog.vl_types.all;
entity Subsystem_tb is
end Subsystem_tb;
